package pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  	`include "transaction.sv"
  	`include "sequence.sv"
  	`include "sequencer.sv"
  	`include "driver.sv"
  	`include "monitor.sv"
	`include "scoreboard.sv";
	`include "coverage.sv"
	`include "agent.sv";
	`include "env.sv";
	`include "base_test.sv"
	`include "apb_read_write_test.sv"
	`include "apb_write_test.sv"
	`include "apb_read_test.sv"
	`include "apb_slverr_test.sv"
    
endpackage

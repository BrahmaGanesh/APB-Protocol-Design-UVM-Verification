class agent extends uvm_agent;
    `uvm_component_utils(agent)

    driver    drv;
    sequencer seqr;
    monitor   mon;

    uvm_active_passive_enum is_active = UVM_ACTIVE;

    function new(string name="agent", uvm_component parent=null);
        super.new(name,parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        mon = monitor::type_id::create("mon", this);

        if (is_active == UVM_ACTIVE) begin
            drv  = driver   ::type_id::create("drv",  this);
            seqr = sequencer::type_id::create("seqr", this);
        end
    endfunction

    function void connect_phase(uvm_phase phase);
        if (is_active == UVM_ACTIVE) begin
        drv.seq_item_port.connect(seqr.seq_item_export);
        end
    endfunction

endclass
